----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:35:50 01/09/2015 
-- Design Name: 
-- Module Name:    logo - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity logo is
    Port ( 
      clk_pixel : IN std_logic;
      --
		i_red     : IN std_logic_vector(7 downto 0);
		i_green   : IN std_logic_vector(7 downto 0);
		i_blue    : IN std_logic_vector(7 downto 0);
		i_blank   : IN std_logic;
		i_hsync   : IN std_logic;
		i_vsync   : IN std_logic;          
      --
		o_red     : OUT std_logic_vector(7 downto 0);
		o_green   : OUT std_logic_vector(7 downto 0);
		o_blue    : OUT std_logic_vector(7 downto 0);
		o_blank   : OUT std_logic;
		o_hsync   : OUT std_logic;
		o_vsync   : OUT std_logic);  
end logo;

architecture Behavioral of logo is

   -------------------------
   -- Part of the pipeline
   -------------------------
	signal a_red     : std_logic_vector(7 downto 0);
	signal a_green   : std_logic_vector(7 downto 0);
	signal a_blue    : std_logic_vector(7 downto 0);
	signal a_blank   : std_logic;
	signal a_hsync   : std_logic;
	signal a_vsync   : std_logic;  

   -------------------------------
   -- Counters for screen position   
   -------------------------------
   signal x : STD_LOGIC_VECTOR (10 downto 0);
   signal y : STD_LOGIC_VECTOR (10 downto 0);

   signal pixel : std_logic_vector(23 downto 0) := (others => '0'); 
   type mem_array is array (0 to 16383) of std_logic_vector(23 downto 0);
   signal address : unsigned(13 downto 0);
   constant logo : mem_array := (
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"818181",x"020202",
x"020202",x"020202",x"020202",x"020202",x"414141",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"818181",x"020202",x"331900",
x"653200",x"653200",x"4c2600",x"000000",x"010101",x"030303",x"030303",x"030303",
x"030303",x"424242",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"818181",x"030303",
x"030303",x"030303",x"030303",x"030303",x"030303",x"020202",x"331900",x"663300",
x"663300",x"663300",x"663300",x"5f2f00",x"201000",x"140a00",x"000000",x"000000",
x"000000",x"010101",x"030303",x"030303",x"030303",x"424242",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"808080",x"000000",
x"321900",x"643200",x"321900",x"000000",x"000000",x"000000",x"010100",x"020100",
x"341a00",x"663300",x"663300",x"2e1700",x"000000",x"04080f",x"172e5b",x"101f3e",
x"000000",x"000000",x"261a0d",x"7c5329",x"714b26",x"010101",x"040404",x"434343",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"828282",x"040404",x"040404",x"040404",x"040404",x"020202",x"000000",
x"331a00",x"663300",x"653300",x"643200",x"643200",x"643200",x"321900",x"000000",
x"010100",x"020100",x"0f0700",x"010000",x"0f1f3c",x"3367cc",x"4080ff",x"2c57ad",
x"101f3e",x"000000",x"000000",x"010100",x"020201",x"000000",x"000000",x"010101",
x"040404",x"040404",x"434343",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"828282",x"030303",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",
x"010100",x"341a00",x"663300",x"663300",x"663300",x"663300",x"331a00",x"000000",
x"000000",x"000000",x"000000",x"0c172d",x"3c77ee",x"4080ff",x"4080ff",x"4080ff",
x"2850a0",x"000000",x"182f5d",x"000000",x"000000",x"282727",x"a19d9d",x"797676",
x"000000",x"000000",x"010101",x"050505",x"050505",x"444444",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"444444",x"050505",x"050505",x"050505",x"050505",
x"030303",x"321900",x"643200",x"643200",x"643200",x"643200",x"643200",x"643200",
x"321900",x"010100",x"020100",x"020100",x"341a00",x"341a00",x"010100",x"504f4f",
x"979494",x"151414",x"000000",x"3467cd",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"1c3971",x"04070f",x"305fbe",x"000000",x"000000",x"706d6d",x"a4a0a0",x"a39f9f",
x"787676",x"000000",x"000000",x"000000",x"000000",x"010101",x"050505",x"050505",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"444444",x"020202",x"000000",x"000000",x"000000",x"000000",
x"000000",x"331a00",x"663300",x"663300",x"663300",x"663300",x"663300",x"663300",
x"331a00",x"000000",x"000000",x"000000",x"010100",x"010100",x"504e4e",x"a29e9e",
x"4a4848",x"000000",x"000000",x"3c78ef",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"0d1932",x"182f5e",x"3060bf",x"000000",x"000000",x"525050",x"a4a0a0",x"a4a0a0",
x"a39f9f",x"787575",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",
x"060606",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"444444",x"020202",x"000000",x"4a2600",x"633200",x"321900",x"000000",
x"000000",x"020100",x"030100",x"351a00",x"663300",x"663300",x"663300",x"351a00",
x"020100",x"504e4e",x"a09c9c",x"a09c9c",x"a09c9c",x"a09c9c",x"a29e9e",x"737070",
x"010101",x"000000",x"13264b",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"1a3366",
x"04070e",x"2f5fbc",x"1d3a73",x"000000",x"000000",x"666363",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a39f9f",x"a09c9c",x"a09c9c",x"a09c9c",x"a09c9c",x"787575",x"000000",
x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"404040",x"000000",x"4a2600",x"653300",x"663300",x"653300",x"633200",
x"633200",x"633200",x"321900",x"020100",x"030100",x"030100",x"351a00",x"331a00",
x"000000",x"525050",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"212020",
x"000000",x"172d5a",x"407ffd",x"4080ff",x"4080ff",x"3971e1",x"162c57",x"000000",
x"1b366c",x"3d79f1",x"050912",x"000000",x"000000",x"8e8b8b",x"a4a0a0",x"807d7d",
x"a4a0a0",x"a4a0a0",x"9b9797",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a39f9f",x"a09c9c",
x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"454545",x"020202",x"4a2600",x"653300",x"663300",x"663300",x"663300",x"663300",
x"663300",x"663300",x"653300",x"321900",x"000000",x"000000",x"020100",x"020100",
x"504e4e",x"a29e9e",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"888585",x"000000",
x"0b162c",x"407ffd",x"4080ff",x"4080ff",x"4080ff",x"407ffd",x"366cd8",x"080f1e",
x"3870df",x"1a3365",x"000000",x"000000",x"000000",x"242323",x"050505",x"000000",
x"050505",x"242323",x"040404",x"2e2d2d",x"888585",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"404040",x"000000",x"4d2600",x"663300",x"663300",x"663300",x"663300",x"663300",
x"663300",x"663300",x"351b00",x"020100",x"504e4e",x"9f9b9b",x"504e4e",x"000000",
x"525050",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"9b9797",x"0d0d0d",x"04070e",
x"376edb",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3f7df9",
x"2c57ad",x"070e1c",x"000000",x"000000",x"000000",x"132549",x"2a54a7",x"172e5c",
x"13264c",x"000000",x"172e5c",x"13264c",x"030303",x"7e7b7b",x"a4a0a0",x"a4a0a0",
x"000000",x"080808",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"464646",x"080808",x"080808",
x"020202",x"000000",x"020200",x"030200",x"030200",x"351b00",x"663300",x"663300",
x"663300",x"351b00",x"020100",x"504e4e",x"a29e9e",x"a4a0a0",x"a29e9e",x"9f9b9b",
x"a29e9e",x"a4a0a0",x"a4a0a0",x"555353",x"050505",x"040404",x"000000",x"1f3e7b",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"3d79f1",x"152a54",x"000000",x"000000",x"1f3d79",x"407ffd",x"4080ff",x"24478d",
x"214182",x"000000",x"204080",x"204080",x"000000",x"141c2a",x"32343b",x"888585",
x"000000",x"000000",x"080808",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"474747",x"020202",x"4a2500",x"623100",
x"623100",x"190c00",x"000000",x"000000",x"000000",x"020100",x"040200",x"351b00",
x"663300",x"331a00",x"4f4d4d",x"a19d9d",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"555353",x"060606",x"030303",x"000000",x"000000",x"04070e",x"386fdd",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3d79f2",
x"162c57",x"000000",x"000000",x"0b162b",x"1d3972",x"4080ff",x"4080ff",x"3163c4",
x"050912",x"000000",x"2f5ebb",x"3467cd",x"000000",x"1c376d",x"102040",x"181717",
x"9e9a9a",x"000000",x"000000",x"090909",x"090909",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"474747",x"4c2702",x"623100",x"653300",x"663300",
x"663300",x"633200",x"623100",x"190c00",x"000000",x"190000",x"190000",x"020100",
x"040200",x"020100",x"525050",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"555353",
x"060606",x"030303",x"0d0d0d",x"0d0d0d",x"000000",x"000000",x"182f5d",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3973e4",x"2a55a9",x"060c17",
x"000000",x"000000",x"000000",x"050b15",x"244890",x"264c97",x"122549",x"010102",
x"000000",x"224386",x"3264c7",x"0a1427",x"04070e",x"3b76eb",x"091122",x"131313",
x"a4a0a0",x"9e9a9a",x"9e9a9a",x"000000",x"000000",x"090909",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"474747",x"030303",x"714b25",x"976431",x"723f0c",x"663300",
x"663300",x"663300",x"663300",x"633200",x"623100",x"321900",x"010000",x"000000",
x"000000",x"000000",x"525050",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"4d4b4b",x"030303",
x"000000",x"000000",x"000000",x"000000",x"0f1e3b",x"000000",x"2b57ad",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"112142",x"000000",x"000000",
x"000000",x"000000",x"000000",x"000000",x"060b15",x"010103",x"000000",x"040810",
x"244890",x"1b356a",x"010103",x"070e1b",x"2e5cb8",x"1e3c77",x"000000",x"767474",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"9e9a9a",x"000000",x"000000",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"404040",x"000000",x"734d26",x"996633",x"986532",x"976431",
x"976431",x"976431",x"723f0c",x"663300",x"1d0e00",x"020100",x"4f4d4d",x"9d9999",
x"9d9999",x"9d9999",x"a19d9d",x"a4a0a0",x"a4a0a0",x"4d4b4b",x"020202",x"000000",
x"000000",x"000000",x"000000",x"000000",x"204080",x"214385",x"3b77ed",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"0c1830",x"000000",x"000000",
x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",
x"000000",x"000000",x"13264b",x"376fdd",x"13254a",x"010103",x"1d1c1c",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"9d9999",x"000000",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"404040",x"000000",x"050302",x"070402",x"754e27",x"996633",
x"996633",x"996633",x"986532",x"976431",x"26190c",x"4f4d4d",x"a19d9d",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"565454",x"020202",x"000000",x"000000",
x"000000",x"000000",x"000000",x"000000",x"23478d",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"040810",x"172d2d",x"7bf4f4",
x"73e4e4",x"5ab4b4",x"4a9494",x"152a2a",x"000000",x"000000",x"000000",x"070f1d",
x"2a54a7",x"204080",x"0a1326",x"020508",x"030303",x"000000",x"292828",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"404040",x"000000",x"492500",x"180c00",x"050402",x"070502",
x"070502",x"070502",x"754e27",x"2c1d0e",x"020101",x"525050",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"353434",x"000000",x"000000",x"000000",
x"070d1a",x"000000",x"000000",x"000000",x"3060bf",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"102040",x"020303",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"7dfafa",x"62c4c4",x"244747",x"000000",x"010203",
x"020508",x"000000",x"101010",x"000000",x"0d0d0d",x"252525",x"020202",x"070707",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"0b0b0b",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"494949",x"030303",x"000000",x"4d2600",x"623200",x"613100",x"613100",
x"180c00",x"000000",x"050402",x"020101",x"000000",x"525050",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"565454",x"020202",x"000000",x"2952a3",x"0b172d",
x"122346",x"000000",x"000000",x"03070d",x"3b77ec",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2b55a9",x"000000",x"6ad2d2",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"7ffcfc",x"4a9393",x"000000",
x"0d0d0d",x"616161",x"656565",x"494949",x"010101",x"0e0e0e",x"252525",x"000000",
x"080808",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"797979",x"131313",x"000000",x"351b00",x"5e2f00",x"663300",x"663300",x"663300",
x"4f2800",x"472400",x"472400",x"120900",x"000000",x"525050",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"6b6868",x"191818",x"000000",x"0f1f3d",x"4080ff",x"050a13",
x"000000",x"000000",x"1b356a",x"366cd6",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3b77ec",x"000000",x"5ab3b3",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"3c7676",
x"000000",x"616161",x"666666",x"5e5e5e",x"353535",x"0d0d0d",x"262626",x"000000",
x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"7a7a7a",
x"131313",x"000000",x"351b00",x"5e2f00",x"663300",x"663300",x"663300",x"663300",
x"663300",x"663300",x"663300",x"1a0d00",x"000000",x"525050",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"6b6868",x"191818",x"000000",x"000000",x"264b95",x"4080ff",x"000000",
x"000000",x"000000",x"1c3870",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"03060d",x"408080",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"7ffcfc",
x"2b5656",x"2a2a2a",x"666666",x"666666",x"4d4d4d",x"040404",x"141414",x"242424",
x"000000",x"313030",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"7a7a7a",x"4d4d4d",x"131313",
x"000000",x"000000",x"4d2600",x"663300",x"663300",x"663300",x"663300",x"663300",
x"663300",x"663300",x"311800",x"080400",x"565353",x"8b8888",x"a4a0a0",x"a4a0a0",
x"6b6969",x"191919",x"181818",x"000000",x"1a3366",x"4080ff",x"356ad3",x"000000",
x"000000",x"000000",x"204080",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3162c3",x"102040",x"408080",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"6edcdc",x"060d0d",x"3d3d3d",x"666666",x"5e5e5e",x"353535",x"0d0d0d",x"333333",
x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"726f6f",x"000000",x"4d4d4d",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"7a7a7a",x"141414",x"351a00",x"472300",
x"472300",x"120900",x"170c00",x"1f1000",x"542a00",x"663300",x"663300",x"663300",
x"311900",x"1f1000",x"080400",x"565353",x"989494",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"525050",x"000000",x"080808",x"000000",x"376edc",x"4080ff",x"3060bf",x"000000",
x"03060c",x"000000",x"3265c8",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"366cd7",x"356ad3",x"264c97",x"102040",x"224343",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"3d7878",x"080808",x"5b5b5b",x"666666",x"4d4d4d",x"040404",x"101010",
x"232323",x"000000",x"323131",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"000000",
x"4e4e4e",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"351a00",x"5e2f00",x"663300",
x"663300",x"4f2700",x"472300",x"120900",x"170c00",x"1f1000",x"1f1000",x"1f1000",
x"080400",x"000000",x"565353",x"989494",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"6b6969",
x"191919",x"242424",x"0d0d0d",x"0b162c",x"4080ff",x"4080ff",x"2d5ab3",x"000000",
x"2a55a8",x"244991",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"3162c3",x"3162c3",x"2f5ebc",x"3366cc",x"1a3568",x"0c1830",x"387070",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"7efcfc",x"0e1c1c",x"363636",x"666666",x"4d4d4d",x"000000",x"000000",
x"333333",x"000000",x"000000",x"323131",x"a4a0a0",x"a4a0a0",x"726f6f",x"726f6f",
x"000000",x"4e4e4e",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"7b7b7b",x"63482e",x"815223",x"6f3c09",x"663300",
x"663300",x"663300",x"663300",x"4e2700",x"462300",x"462300",x"120900",x"000000",
x"555353",x"716f6f",x"979494",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"525050",
x"232323",x"565656",x"000000",x"1e3c78",x"356ad3",x"4080ff",x"3366cc",x"0b162c",
x"254a93",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3972e3",x"3870df",
x"3972e3",x"3060bf",x"3060bf",x"3060bf",x"3d7af3",x"3060bf",x"13264c",x"204040",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"346868",x"020202",x"666666",x"5e5e5e",x"353535",x"000000",
x"333333",x"232323",x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"404040",x"24180c",x"7f552a",x"8d5a27",x"895623",
x"895623",x"6f3c09",x"663300",x"663300",x"663300",x"321900",x"080400",x"555353",
x"979494",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"6c6969",x"1a1919",
x"333333",x"434343",x"000000",x"3366cb",x"3468cf",x"4080ff",x"3f7efb",x"1f3e7c",
x"274e9c",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3366cb",x"2d5ab3",
x"3060bf",x"24488f",x"3060bf",x"3c78ef",x"3060bf",x"2c58af",x"1c3870",x"204040",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"7efbfb",x"1c3838",x"3d3d3d",x"666666",x"4d4d4d",x"000000",
x"101010",x"333333",x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"716e6e",x"000000",x"4f4f4f",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"c3c3c3",x"2c2c2c",x"24180c",x"7f552a",x"996633",
x"996633",x"8d5a27",x"895623",x"895623",x"895623",x"221609",x"000000",x"7b7878",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"6c6969",x"1a1919",x"232323",
x"565656",x"1b1b1b",x"0b162c",x"4080ff",x"3060bf",x"4080ff",x"4080ff",x"274e9b",
x"214284",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2c58af",
x"3060bf",x"3870df",x"2d5ab4",x"2952a4",x"2952a4",x"3b76eb",x"112244",x"204040",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"56abab",x"1d1d1d",x"666666",x"4d4d4d",x"000000",
x"000000",x"333333",x"232323",x"000000",x"333232",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"000000",x"24180c",x"302010",
x"302010",x"302010",x"7f552a",x"996633",x"996633",x"261a0d",x"000000",x"7b7878",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"525050",x"000000",x"333333",
x"666666",x"080808",x"102040",x"4080ff",x"3f7efb",x"4080ff",x"4080ff",x"3b76eb",
x"366cd7",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2f5ebb",
x"3b76eb",x"3366cb",x"23468b",x"244890",x"23468b",x"4080ff",x"091224",x"204040",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"7efbfb",x"0e1c1c",x"4a4a4a",x"5e5e5e",x"464646",
x"000000",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"351a00",x"462300",x"462300",
x"120900",x"000000",x"24180c",x"302010",x"302010",x"0c0804",x"000000",x"7b7878",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"504e4e",x"1a1a1a",x"232323",x"565656",
x"4a4a4a",x"000000",x"1a3467",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"3b76eb",x"2a54a7",x"3b76eb",x"3972e4",x"000000",x"2e5b5b",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"3c7777",x"282828",x"666666",x"666666",
x"000000",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"190c00",x"552a00",x"663300",
x"4d2700",x"452300",x"452300",x"110900",x"000000",x"000000",x"000000",x"7b7878",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"292828",x"000000",x"333333",x"666666",
x"333333",x"000000",x"2c58af",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"214284",x"000000",x"3a7474",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"6edbdb",x"1a1a1a",x"666666",x"666666",
x"000000",x"101010",x"333333",x"232323",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"341a00",x"5e2f00",x"663300",
x"663300",x"663300",x"663300",x"4d2700",x"452300",x"110900",x"000000",x"7b7878",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"292828",x"232323",x"565656",x"666666",
x"333333",x"0b162b",x"3060bf",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"376dd9",x"070d19",x"000000",x"448686",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"203d3d",x"666666",x"666666",
x"000000",x"000000",x"333333",x"333333",x"000000",x"353333",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"adadad",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"7d7d7d",x"151515",x"4d2600",x"663300",x"663300",
x"663300",x"663300",x"663300",x"663300",x"663300",x"1a0d00",x"000000",x"7b7878",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"514f4f",x"0d0d0d",x"333333",x"666666",x"666666",
x"333333",x"102040",x"254a94",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"152a54",x"000000",x"000000",x"6edbdb",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"448686",x"4e4e4e",x"666666",
x"000000",x"000000",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"404040",x"341a00",x"5e2f00",x"663300",x"663300",
x"663300",x"663300",x"663300",x"663300",x"663300",x"1a0d00",x"000000",x"7b7878",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"292828",x"000000",x"333333",x"666666",x"666666",
x"333333",x"183060",x"204080",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"20407e",x"010305",x"000000",x"000000",x"65c9c9",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"66caca",x"2a2a2a",x"666666",
x"000000",x"000000",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"535353",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"7e7e7e",x"535353",x"151515",x"190d00",x"211100",x"211100",x"211100",
x"552b00",x"663300",x"663300",x"663300",x"663300",x"1a0d00",x"535151",x"979393",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"292828",x"343434",x"565656",x"666666",x"666666",
x"333333",x"102040",x"3263c6",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"102040",x"000000",x"000000",x"000000",x"1d3a3a",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"73e4e4",x"020202",x"5b5b5b",
x"000000",x"000000",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"7f7f7f",x"151515",x"331a00",x"442200",x"442200",x"442200",x"442200",x"110900",
x"1a0d00",x"221100",x"221100",x"552b00",x"331a00",x"090400",x"7b7878",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"525050",x"0e0d0d",x"4d4d4d",x"666666",x"666666",x"666666",
x"333333",x"183060",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"102040",x"000000",x"000000",x"000000",x"000000",
x"7bf4f4",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"6edada",x"060b0b",x"353535",
x"444444",x"000000",x"333333",x"333333",x"222222",x"000000",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"6e6b6b",x"000000",x"545454",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"404040",x"331a00",x"5e2f00",x"663300",x"663300",x"663300",x"663300",x"4d2600",
x"442200",x"442200",x"442200",x"2b1500",x"090400",x"535050",x"979393",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"292828",x"000000",x"4d4d4d",x"666666",x"666666",x"666666",
x"333333",x"102040",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"2851a0",x"0f1e3b",x"23468b",x"03060b",x"000000",
x"60bfbf",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"3e7b7b",x"333333",
x"666666",x"000000",x"333333",x"333333",x"333333",x"000000",x"363535",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"404040",x"66401a",x"6f3c09",x"663300",x"663300",x"663300",x"663300",x"663300",
x"663300",x"663300",x"331a00",x"090400",x"525050",x"969393",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"292828",x"333333",x"5e5e5e",x"666666",x"666666",x"666666",
x"333333",x"102040",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"13254a",x"000000",
x"56aaaa",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"3d7a7a",x"0b0b0b",
x"555555",x"000000",x"333333",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"404040",x"261a0d",x"73481e",x"885522",x"885522",x"6f3c09",x"663300",x"663300",
x"663300",x"663300",x"1a0d00",x"525050",x"969393",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"525151",x"0e0e0e",x"4d4d4d",x"666666",x"666666",x"666666",x"666666",
x"404040",x"0d1b35",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2f5dba",x"000000",
x"204040",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"509f9f",x"000000",
x"4d4d4d",x"000000",x"333333",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"404040",x"000000",x"261a0d",x"80552b",x"996633",x"8c5926",x"885522",x"885522",
x"885522",x"3c2209",x"5a5450",x"969393",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"292828",x"000000",x"4d4d4d",x"666666",x"666666",x"666666",x"666666",
x"4a4a4a",x"000000",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"376dda",x"000000",
x"3d7a7a",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"60bfbf",x"000000",
x"1a1a1a",x"000000",x"333333",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",
x"a4a0a0",x"373636",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"8f8f8f",x"1a1a1a",x"000000",x"442d17",x"5a3c1e",x"5a3c1e",x"5a3c1e",x"895c2e",
x"996633",x"261a0d",x"494747",x"939090",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"292828",x"000000",x"4d4d4d",x"666666",x"666666",x"666666",x"666666",
x"4d4d4d",x"000000",x"366bd5",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"172d5a",
x"408080",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"60bfbf",x"000000",
x"000000",x"000000",x"333333",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"696969",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"404040",x"000000",x"201000",x"2a1500",x"2a1500",x"2a1500",x"4e3217",
x"5a3c1e",x"170f08",x"000000",x"7b7878",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"292828",x"000000",x"4d4d4d",x"666666",x"666666",x"666666",x"666666",
x"4d4d4d",x"000000",x"3060bf",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"376edb",x"2e5cb7",x"3971e1",x"366cd7",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"1f3d7a",
x"2e5c5c",x"54a7a7",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"6dd9d9",x"000000",
x"000000",x"000000",x"333333",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",
x"615f5f",x"000000",x"686868",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"404040",x"000000",x"4d2600",x"663300",x"663300",x"663300",x"391d00",
x"2a1500",x"2a1500",x"0b0500",x"494747",x"939090",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"292828",x"000000",x"4d4d4d",x"666666",x"666666",x"666666",x"666666",
x"5d5d5d",x"000000",x"264b95",x"3263c5",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"3e7bf5",x"0b162c",x"000000",x"020306",x"000000",
x"0a1427",x"1e3c77",x"3161c1",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"204080",
x"000000",x"0d1a1a",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"6bd5d5",x"000000",
x"000000",x"000000",x"333333",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",
x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"404040",x"000000",x"4d2600",x"663300",x"663300",x"663300",x"663300",
x"663300",x"663300",x"381d00",x"0a0500",x"4a4747",x"949090",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"292828",x"000000",x"4d4d4d",x"666666",x"666666",x"666666",x"666666",
x"4f4f4f",x"000000",x"204080",x"376dd9",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"2c58af",x"000000",x"000000",x"000000",x"040810",
x"0c172d",x"000000",x"060b16",x"376edc",x"4080ff",x"4080ff",x"4080ff",x"3162c3",
x"0d1a34",x"204040",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"6dd9d9",x"000000",
x"000000",x"000000",x"333333",x"333333",x"333333",x"000000",x"424141",x"a4a0a0",
x"000000",x"676767",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"b2b2b2",x"262626",x"000000",x"4d2600",x"663300",x"663300",x"663300",x"663300",
x"663300",x"663300",x"663300",x"381d00",x"0a0500",x"7b7878",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"292828",x"101010",x"525252",x"666666",x"666666",x"666666",x"666666",
x"4d4d4d",x"000000",x"1c3870",x"3a73e5",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"24488f",x"000000",x"284f9d",x"224487",x"000000",
x"3468cf",x"14274d",x"000000",x"070e1c",x"376edc",x"4080ff",x"4080ff",x"4080ff",
x"162b56",x"336666",x"5cb8b8",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"000000",
x"000000",x"000000",x"333333",x"333333",x"1e1e1e",x"000000",x"a4a0a0",x"a4a0a0",
x"000000",x"989898",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"b3b3b3",
x"262626",x"2e1f0f",x"3d2914",x"3d2205",x"3d1f00",x"3d1f00",x"3d1f00",x"3d1f00",
x"5c2e00",x"663300",x"663300",x"472400",x"413830",x"8c8888",x"a4a0a0",x"a4a0a0",
x"737070",x"191818",x"262626",x"595959",x"666666",x"666666",x"666666",x"666666",
x"4d4d4d",x"000000",x"162b56",x"3060bf",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"376dd9",x"000000",x"264b96",x"4080ff",x"203f7d",
x"1b376c",x"3b75e9",x"03050a",x"000000",x"13274d",x"4080ff",x"4080ff",x"4080ff",
x"0e1b36",x"000000",x"000000",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"78efef",x"000000",
x"000000",x"000000",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",x"a4a0a0",
x"424040",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"6e5f4f",
x"3d2914",x"82572b",x"996633",x"54381c",x"3d2914",x"0f0a05",x"000000",x"000000",
x"2e1700",x"5c2e00",x"472400",x"0f0800",x"7b7878",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"292828",x"000000",x"262626",x"595959",x"666666",x"666666",x"666666",x"666666",
x"3c3c3c",x"000000",x"142850",x"3f7df9",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"070d1a",x"0b172d",x"4080ff",x"376dd9",
x"020306",x"4080ff",x"254a93",x"070d1a",x"070d1a",x"3367cc",x"4080ff",x"3367cc",
x"000000",x"000000",x"000000",x"7bf6f6",x"6ad3d3",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"78efef",x"000000",
x"000000",x"141414",x"333333",x"333333",x"000000",x"000000",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"999999",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"c29b75",
x"9e6b38",x"996633",x"996633",x"996633",x"996633",x"54381c",x"3d2914",x"3d2914",
x"0f0a05",x"4d2600",x"1a0d00",x"313030",x"8b8888",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"292828",x"000000",x"262626",x"595959",x"666666",x"666666",x"666666",x"666666",
x"2d2d2d",x"050a13",x"1f3e7c",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"1d3a72",x"000000",x"2c57ad",x"4080ff",
x"193365",x"4080ff",x"3a75e9",x"172e5c",x"1a3569",x"1e3b76",x"4080ff",x"204080",
x"020509",x"1d3b75",x"020509",x"274d4d",x"132727",x"80ffff",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"78efef",x"000000",
x"000000",x"292929",x"313131",x"1f1f1f",x"000000",x"414040",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"9c856e",
x"a17345",x"ad7a47",x"ad7a47",x"ad7a47",x"9e6b38",x"996633",x"996633",x"996633",
x"54381c",x"3e2105",x"40372f",x"8b8888",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"292828",x"000000",x"262626",x"595959",x"666666",x"666666",x"666666",x"666666",
x"373737",x"204080",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3a75e9",x"020509",x"080f1d",x"386fdd",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3265c9",x"060b17",x"4080ff",x"3d7af2",
x"3366cc",x"4080ff",x"102040",x"030707",x"000000",x"7bf6f6",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"000000",
x"050a13",x"050a13",x"090d16",x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",
x"5d462f",x"7c5d3e",x"b88a5c",x"cc9966",x"b5824f",x"ad7a47",x"ad7a47",x"9e6b38",
x"996633",x"261a0d",x"7b7878",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"292828",x"000000",x"262626",x"595959",x"666666",x"666666",x"666666",x"666666",
x"4d4d4d",x"122447",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"214182",x"000000",x"162c57",
x"4080ff",x"4080ff",x"3a74e6",x"3c77ed",x"1d3b74",x"000000",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"1e3d79",x"000000",x"000000",x"60bfbf",x"80ffff",x"80ffff",
x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"000000",
x"204080",x"204080",x"3a75e9",x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"8b8b8b",
x"646464",x"191919",x"5d462f",x"7c5d3e",x"7c5d3e",x"7c5d3e",x"b88a5c",x"b5824f",
x"ad7a47",x"2b1f12",x"7b7878",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"292828",x"000000",x"262626",x"4a4a4a",x"616161",x"666666",x"666666",x"666666",
x"575757",x"020407",x"3a74e6",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3a75e8",x"060d19",x"102040",
x"4080ff",x"4080ff",x"366dd8",x"183060",x"000000",x"0d1932",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"224589",x"020509",x"0a1529",x"448686",x"80ffff",x"80ffff",
x"6fdddd",x"6fdddd",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"000000",
x"1e3c77",x"122447",x"284f9d",x"000000",x"403f3f",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"646161",x"000000",x"646464",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"8a8a8a",x"191919",x"000000",x"000000",x"000000",x"5e462f",x"7d5d3e",
x"b88a5c",x"33261a",x"4b4a4a",x"949191",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"292828",x"000000",x"171717",x"2e2e2e",x"595959",x"666666",x"666666",x"666666",
x"666666",x"0a0a0a",x"182f5e",x"4080ff",x"4080ff",x"4080ff",x"3a74e6",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"102040",x"0a1427",
x"4080ff",x"3c78ef",x"3870df",x"1e3c77",x"000000",x"204080",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"3a75e8",x"23468a",x"102040",x"408080",x"80ffff",x"80ffff",
x"244747",x"346767",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"000000",
x"1e3d79",x"224589",x"060c17",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"646262",
x"000000",x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"404040",x"000000",x"1e0f00",x"281400",x"281400",x"281400",
x"684c2f",x"1f1810",x"000000",x"4b4a4a",x"949191",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"595757",x"101010",x"000000",x"262626",x"595959",x"666666",x"666666",x"666666",
x"666666",x"1a1a1a",x"254991",x"4080ff",x"4080ff",x"4080ff",x"3e7df8",x"3e7cf6",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"102040",x"000000",
x"4080ff",x"3e7cf6",x"366cd6",x"1e3d79",x"000000",x"204080",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"0a1529",x"387070",x"80ffff",x"80ffff",
x"2d5959",x"1c3737",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"80ffff",x"000000",
x"1e3c77",x"0c172e",x"000000",x"403e3e",x"a4a0a0",x"a4a0a0",x"646262",x"000000",
x"636363",x"636363",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"898989",x"191919",x"4d2600",x"663300",x"663300",x"663300",
x"371c00",x"271400",x"271400",x"0a0500",x"4c4a4a",x"949191",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"292828",x"000000",x"262626",x"595959",x"666666",x"666666",x"666666",
x"666666",x"1a1a1a",x"224487",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3e7df8",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"102040",x"000000",
x"4080ff",x"3060bf",x"3468cf",x"204080",x"000000",x"224488",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"08101f",x"408080",x"57adad",x"63c6c6",
x"408080",x"000000",x"7cf7f7",x"80ffff",x"80ffff",x"80ffff",x"74e7e7",x"000000",
x"020407",x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"656262",x"000000",x"626262",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"404040",x"4d2600",x"663300",x"663300",x"663300",
x"663300",x"663300",x"663300",x"371c00",x"0a0500",x"4c4a4a",x"949191",x"a4a0a0",
x"a4a0a0",x"292828",x"000000",x"262626",x"595959",x"666666",x"666666",x"666666",
x"666666",x"3a3a3a",x"0c182f",x"4080ff",x"3c78ef",x"3a74e7",x"3870df",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"102040",x"000000",
x"4080ff",x"3e7cf8",x"2c58af",x"204080",x"000000",x"3060bf",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"3a74e7",x"000000",x"448888",x"081010",x"040707",
x"61c1c1",x"000000",x"60bfbf",x"80ffff",x"80ffff",x"80ffff",x"60bfbf",x"000000",
x"000000",x"000000",x"3f3d3d",x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"b6b6b6",x"282828",x"4d2600",x"663300",x"663300",x"663300",
x"663300",x"663300",x"663300",x"663300",x"371b00",x"0a0500",x"7b7878",x"a4a0a0",
x"a4a0a0",x"585656",x"100f0f",x"181818",x"464646",x"5d5d5d",x"666666",x"666666",
x"666666",x"636363",x"0d0d0d",x"2a53a6",x"4080ff",x"3870df",x"3a74e7",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"1a3468",x"000000",
x"4080ff",x"4080ff",x"3468cf",x"1c3870",x"000000",x"3a74e8",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"224487",x"000000",x"234747",x"000000",x"000000",
x"64c7c7",x"040808",x"4c9797",x"80ffff",x"80ffff",x"80ffff",x"4c9797",x"000000",
x"000000",x"000000",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"b6b6b6",x"282828",x"000000",x"2f1800",x"3f2000",x"5c2e00",x"663300",
x"663300",x"663300",x"663300",x"663300",x"663300",x"1a0d00",x"7b7878",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"292828",x"000000",x"262626",x"434343",x"5d5d5d",x"666666",
x"666666",x"666666",x"464646",x"060c18",x"3060bf",x"3060bf",x"3a74e8",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"264c98",x"000000",
x"4080ff",x"3e7cf7",x"3a74e8",x"183060",x"000000",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"224488",x"000000",x"000000",x"060c18",x"000000",
x"1b3737",x"0c1818",x"182f2f",x"407f7f",x"68cfcf",x"78efef",x"1c3737",x"000000",
x"000000",x"3e3d3d",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"b7b7b7",x"282828",x"2c1d0e",x"3a2713",x"3a2713",x"0f0a05",x"2f1800",x"3f2000",
x"3f2000",x"5c2e00",x"663300",x"663300",x"663300",x"1a0d00",x"7b7878",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"292828",x"000000",x"262626",x"333333",x"4d4d4d",x"666666",
x"666666",x"666666",x"5c5c5c",x"000000",x"081020",x"2a54a7",x"3a74e7",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3264c7",x"000000",
x"3a74e7",x"3e7cf7",x"3e7cf7",x"204080",x"060c18",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"366cd7",x"040810",x"2850a0",x"204080",x"000000",
x"040808",x"346868",x"000000",x"5cb8b8",x"80ffff",x"80ffff",x"204040",x"000000",
x"3e3c3c",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"404040",x"2c1d0e",x"81562b",x"996633",x"996633",x"52361b",x"3a2613",x"3a2613",
x"0f0a05",x"301800",x"402000",x"402000",x"402000",x"100800",x"7b7878",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"292828",x"000000",x"262626",x"333333",x"434343",x"5d5d5d",
x"666666",x"666666",x"636363",x"000000",x"000000",x"224488",x"2c58af",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"020408",
x"3468cf",x"4080ff",x"3468cf",x"204080",x"102040",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3870e0",x"4080ff",x"3e7cf7",x"142850",
x"040808",x"78efef",x"000000",x"4c9797",x"78efef",x"509f9f",x"142828",x"000000",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"000000",x"000000",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"404040",x"654322",x"86592d",x"996736",x"9f6c39",x"9b6835",x"996633",x"996633",
x"352311",x"130d06",x"130d06",x"130d06",x"050302",x"0f0f0f",x"807d7d",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"383737",x"050505",x"222222",x"303030",x"333333",x"4a4a4a",
x"636363",x"666666",x"666666",x"131313",x"000000",x"102040",x"3e7cf7",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"264c97",
x"3a74e7",x"4080ff",x"366cd7",x"264c97",x"102040",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3264c7",
x"000000",x"54a8a8",x"204040",x"285050",x"204040",x"000000",x"000000",x"000000",
x"716e6e",x"908c8c",x"a4a0a0",x"a4a0a0",x"908c8c",x"000000",x"181818",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"575757",x"080808",x"000000",x"866544",x"c69463",x"aa7744",x"9f6c39",x"9f6c39",
x"9f6c39",x"9b6835",x"996633",x"8b5d2f",x"31251a",x"807d7d",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"292828",x"000000",x"1a1a1a",x"333333",x"333333",
x"4d4d4d",x"666666",x"666666",x"434343",x"040810",x"2c58af",x"3c78ef",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"366cd7",x"1e3c77",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3e7cf7",
x"0c1830",x"285050",x"306060",x"000000",x"1e3c77",x"3870df",x"3060bf",x"18305f",
x"040810",x"000000",x"343232",x"908d8d",x"000000",x"000000",x"474747",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"575757",x"1f1f1f",x"080808",x"876544",x"b4875a",x"b4875a",x"c69563",
x"cc9966",x"aa7744",x"9f6c39",x"281b0e",x"7b7878",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"292828",x"000000",x"171717",x"303030",x"333333",
x"4a4a4a",x"606060",x"636363",x"636363",x"0a0a0a",x"244990",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"2c58af",x"000000",x"000000",x"000000",x"0e1d39",x"2851a1",x"142951",x"142951",
x"102141",x"000000",x"000000",x"000000",x"000000",x"1f1f1f",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"565656",x"1e1e1e",x"080808",x"000000",x"876544",
x"b4875a",x"b4875a",x"c69563",x"453423",x"736e6d",x"9f9b9b",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"373636",x"050505",x"000000",x"1a1a1a",x"333333",
x"333333",x"333333",x"4a4a4a",x"636363",x"333333",x"060c18",x"3a74e8",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3c79f0",
x"183161",x"000000",x"000000",x"000000",x"000000",x"04080f",x"14274e",x"182f5e",
x"1c376e",x"182f5e",x"0c172e",x"020408",x"000000",x"919191",x"f8f8f8",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"000000",x"120e09",
x"060503",x"000000",x"876544",x"b4875a",x"2d2217",x"6d6a6a",x"9f9b9b",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"373636",x"0a0a0a",x"171717",x"303030",
x"333333",x"333333",x"333333",x"4a4a4a",x"595959",x"131313",x"172d59",x"3e7cf8",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3a74e8",x"091121",
x"000000",x"020408",x"04080f",x"102040",x"23478d",x"102040",x"3e7cf8",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"3a73e6",x"1b376d",x"020408",x"3a3a3a",x"e8e8e8",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"000000",x"99734d",
x"443323",x"17110c",x"060403",x"000000",x"000000",x"000000",x"6d6b6b",x"918e8e",
x"918e8e",x"918e8e",x"9f9c9c",x"a4a0a0",x"a4a0a0",x"5c5959",x"0a0909",x"171717",
x"303030",x"333333",x"333333",x"333333",x"4a4a4a",x"3c3c3c",x"000000",x"264c98",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"172d5a",x"000000",
x"172f5d",x"3973e6",x"3468ce",x"020407",x"3870df",x"3870de",x"3264c7",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2d5bb6",x"020407",x"2a2a2a",
x"d9d9d9",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"000000",x"99734d",
x"cc9966",x"cc9966",x"443322",x"17110b",x"17110b",x"17110b",x"17110b",x"060403",
x"000000",x"000000",x"7b7878",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"525050",x"000000",
x"1a1a1a",x"333333",x"333333",x"333333",x"333333",x"4a4a4a",x"101010",x"0d1932",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2951a1",x"000000",x"274f9c",
x"4080ff",x"4080ff",x"4080ff",x"356bd5",x"3870df",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"214283",x"020509",x"000000",
x"090909",x"c8c8c8",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"555555",x"070707",x"9e7b55",
x"d2a471",x"d2a471",x"ce9c69",x"cc9966",x"cc9966",x"cc9966",x"cc9966",x"443322",
x"16110b",x"060403",x"6e6b6b",x"a09c9c",x"a4a0a0",x"a4a0a0",x"5b5959",x"090909",
x"171717",x"303030",x"333333",x"333333",x"333333",x"333333",x"262626",x"000000",
x"3161c1",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"3972e3",x"2d5ab3",x"0d1932",x"193365",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3e7df8",x"3569d1",x"4080ff",
x"4080ff",x"4080ff",x"3e7df8",x"3162c3",x"193263",x"070707",x"000000",x"000000",
x"000000",x"3a3a3a",x"e1e1e1",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"aaaa89",
x"f8f8c7",x"ffffcc",x"ddbb88",x"d2a471",x"ce9c69",x"cc9966",x"cc9966",x"cc9966",
x"cc9966",x"443322",x"060403",x"6e6b6b",x"a09c9c",x"a4a0a0",x"a4a0a0",x"5b5959",
x"090909",x"171717",x"303030",x"333333",x"333333",x"333333",x"333333",x"050505",
x"0d1932",x"4080ff",x"4080ff",x"4080ff",x"2a55a8",x"3c78ef",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"172e5c",x"000000",x"000000",x"2951a2",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"376eda",x"3e7df8",x"3e7cf6",x"1c376e",x"4080ff",
x"4080ff",x"4080ff",x"193162",x"000000",x"000000",x"505050",x"101010",x"000000",
x"000000",x"000000",x"808080",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"545454",x"070707",
x"abab89",x"e4e4b6",x"e4e4b6",x"f8f8c7",x"ddbb88",x"d1a471",x"d1a471",x"cd9c69",
x"cc9966",x"cc9966",x"33261a",x"000000",x"7b7878",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"5b5959",x"090909",x"171717",x"313131",x"333333",x"333333",x"333333",x"212121",
x"000000",x"3161c2",x"4080ff",x"3265c8",x"3060bf",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"172e5b",x"020407",x"020509",x"2952a4",
x"4080ff",x"4080ff",x"4080ff",x"214384",x"2a54a6",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"102040",x"000000",x"000000",x"696969",x"101010",x"000000",
x"000000",x"000000",x"808080",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"545454",
x"070707",x"000000",x"000000",x"abab89",x"e4e4b7",x"e4e4b7",x"f8f8c7",x"ddbb88",
x"d1a471",x"cd9c69",x"33261a",x"000000",x"7b7878",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"5b5959",x"090909",x"171717",x"2e2e2e",x"2e2e2e",x"313131",x"333333",
x"080808",x"091223",x"366dd9",x"3060bf",x"3263c6",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3162c3",x"13254a",x"000000",
x"2e5db9",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"214284",x"000000",x"000000",x"000000",x"000000",x"000000",
x"04070e",x"060b17",x"696969",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"535353",x"1a1a1a",x"1a1a1a",x"070707",x"000000",x"000000",x"acac89",x"e5e5b7",
x"e5e5b7",x"d6b482",x"34291c",x"0d0c0c",x"7f7c7c",x"a4a0a0",x"a4a0a0",x"a4a0a0",
x"a4a0a0",x"a4a0a0",x"5b5858",x"090808",x"000000",x"000000",x"171717",x"2e2e2e",
x"0c0c0c",x"000000",x"2a55a9",x"2c58af",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2b55aa",
x"3a73e6",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"376dda",x"2b55aa",x"274d9a",x"274d9a",x"3365ca",
x"386fdd",x"0e1d39",x"767676",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"535353",x"1a1a1a",x"070707",x"000000",x"000000",
x"000000",x"acac8a",x"39392e",x"6f6c6c",x"949090",x"949090",x"949090",x"949090",
x"9c9898",x"a4a0a0",x"a4a0a0",x"5a5858",x"101010",x"080808",x"000000",x"000000",
x"000000",x"122346",x"204080",x"366bd6",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"000000",x"808080",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"404040",x"000000",x"0f0b08",
x"140f0a",x"050403",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",
x"525050",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"5a5858",x"101010",x"080808",
x"000000",x"03050a",x"264b96",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"000000",x"a6a6a6",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"535353",x"060606",x"9d7a54",
x"d1a370",x"473c2b",x"15120d",x"140f0a",x"140f0a",x"140f0a",x"140f0a",x"0a0805",
x"4a4949",x"9c9999",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"565454",
x"000000",x"172e5c",x"3a73e5",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3f7df9",x"366cd6",
x"2a54a7",x"2a54a7",x"2a54a7",x"3a74e6",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"376dd9",x"000000",x"bfbfbf",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"525252",x"b3b391",
x"e7e7b9",x"f9f9c7",x"ddba87",x"d1a370",x"d1a370",x"d1a370",x"cf9e6b",x"664d33",
x"000000",x"525050",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"a4a0a0",x"949090",
x"000000",x"1b356a",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2e5cb7",x"0c172d",x"000000",
x"000000",x"000000",x"000000",x"000000",x"1a3467",x"3b75e9",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"274d99",x"000000",x"c5c5c5",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"525252",
x"181818",x"b3b391",x"e7e7b9",x"e7e7b9",x"e7e7b9",x"f3f3c3",x"e8d19e",x"755d41",
x"0c0c0a",x"525050",x"a4a0a0",x"a4a0a0",x"9d9999",x"959191",x"959191",x"9d9999",
x"3f3d3d",x"03050a",x"376dd9",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2d5ab4",x"000000",x"000000",x"000000",
x"000000",x"000000",x"000000",x"000000",x"000000",x"2c58af",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"1b356a",x"363636",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"515151",x"171717",x"171717",x"060606",x"74745d",x"e8e8ba",x"e8e8ba",
x"74745d",x"4b4949",x"959292",x"959292",x"4b4949",x"000000",x"000000",x"4b4949",
x"8c8989",x"0e0e0e",x"214284",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"0d1a34",x"000000",x"000000",x"000000",
x"000000",x"000000",x"000000",x"000000",x"060b16",x"3a73e5",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"0b152a",x"8b8b8b",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"515151",x"171717",x"171717",x"0c0c0c",
x"000000",x"000000",x"000000",x"000000",x"000000",x"0c0c09",x"0c0c09",x"000000",
x"525050",x"414040",x"0b152a",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"000000",x"000000",x"000000",x"000000",
x"161616",x"c6c6c6",x"616161",x"000000",x"254991",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3b75ea",
x"000000",x"d5d5d5",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"8b8b8b",
x"161616",x"161616",x"161616",x"161616",x"0b0b0b",x"75755d",x"75755d",x"000000",
x"4b4949",x"858282",x"070707",x"2d5bb4",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"000000",x"000000",x"000000",x"000000",
x"3a3a3a",x"f4f4f4",x"4f4f4f",x"1e3b76",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"214384",
x"000000",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"808080",x"000000",x"000000",x"000000",
x"000000",x"525050",x"525050",x"0e1b35",x"3f7dfa",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"112346",x"040811",x"000000",x"000000",
x"010306",x"1e283a",x"244890",x"366bd5",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"0b152b",
x"2b2b2b",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"eaeaea",x"d5d5d5",x"6b6b6b",x"000000",
x"000000",x"0e0e0e",x"0e0e0e",x"000000",x"264b95",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"1c386f",x"3d7bf5",x"254b95",x"152b55",
x"2f5eba",x"3e7bf5",x"244890",x"3366ca",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3f7dfa",x"000000",
x"858585",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"eaeaea",x"d4d4d4",
x"d4d4d4",x"d4d4d4",x"d4d4d4",x"848484",x"070e1b",x"3a73e5",x"4080ff",x"4080ff",
x"4080ff",x"366bd5",x"3a73e5",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3468cf",x"2851a0",x"2c59b0",x"091325",
x"274e9a",x"274e9a",x"2952a4",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"142950",x"3a3a3a",
x"f4f4f4",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"2a2a2a",x"122346",x"3f7efa",x"4080ff",
x"4080ff",x"0e1b36",x"2d5bb5",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3f7efa",x"3365ca",x"0d1b35",x"2b55aa",
x"2b55aa",x"24488f",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"2c59b0",x"000000",x"959595",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"d9d9d9",x"151515",x"1c3971",x"3366cc",
x"2e5bb6",x"000000",x"264b96",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"366bd5",x"3d7bf4",x"274e9b",x"2b55a9",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3061c1",x"03060b",x"000000",x"d4d4d4",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"7e7e7e",x"000000",x"000000",
x"0e1b36",x"000000",x"28509e",x"4080ff",x"4080ff",x"3e7bf6",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"274d99",x"4080ff",x"274d99",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"081020",x"000000",x"353535",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"626262",x"000000",
x"000000",x"172d59",x"4080ff",x"4080ff",x"2c58af",x"0a1427",x"3a74e6",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"13264b",x"000000",x"646464",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"5e5e5e",
x"000000",x"2d5ab4",x"4080ff",x"4080ff",x"4080ff",x"0d1a35",x"060c17",x"3a74e6",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"3f7efb",x"000000",x"000000",x"848484",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"bfbfbf",
x"000000",x"3060bf",x"4080ff",x"4080ff",x"4080ff",x"112244",x"000000",x"060c17",
x"305fbe",x"3e7cf6",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"264c97",x"000000",x"000000",x"bfbfbf",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"bfbfbf",
x"000000",x"3d7af4",x"4080ff",x"4080ff",x"4080ff",x"23468b",x"040810",x"000000",
x"000000",x"0f1e3b",x"4080ff",x"4080ff",x"3c77ee",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"3b76eb",x"070e1c",x"010204",x"010204",x"bfbfbf",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"bfbfbf",
x"000000",x"4080ff",x"4080ff",x"4080ff",x"3162c3",x"0b162c",x"000000",x"000000",
x"000000",x"1a3468",x"4080ff",x"1d3a73",x"050a14",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"3f7efb",x"112243",x"010204",x"274e9c",x"102040",x"c4c4c4",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"bfbfbf",
x"000000",x"376edb",x"4080ff",x"3b76eb",x"172e5c",x"112244",x"081020",x"000000",
x"010204",x"356ad3",x"3b76eb",x"03060c",x"224488",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",
x"3a74e7",x"152a53",x"050a14",x"193264",x"4080ff",x"102040",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"bfbfbf",
x"000000",x"1d3a74",x"3c78ef",x"152a54",x"23468b",x"040810",x"000000",x"000000",
x"1f3e7b",x"4080ff",x"152a54",x"091224",x"3d7af3",x"4080ff",x"4080ff",x"4080ff",
x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"4080ff",x"3468d0",x"204080",
x"060c18",x"050a14",x"1d3a74",x"172e5c",x"4080ff",x"03060c",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"e3e3e3",
x"000000",x"000000",x"183060",x"040810",x"091224",x"0b162c",x"020408",x"1c386f",
x"4080ff",x"2c58b0",x"000000",x"03060c",x"0c1830",x"142850",x"204080",x"2c58b0",
x"2c58b0",x"3060c0",x"2c58b0",x"2c58b0",x"244890",x"0c1830",x"000000",x"000000",
x"181c24",x"274e9b",x"3264c7",x"214284",x"3b76eb",x"202020",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"5b5b5b",x"000000",x"142850",x"2c58b0",x"2c58ae",x"2c58ae",x"366cd7",x"3973e4",
x"183161",x"040404",x"6e6e6e",x"7e7e7e",x"5e5e5e",x"2f2f2f",x"0f0f0f",x"0f0f0f",
x"080808",x"040404",x"0f0f0f",x"000000",x"0f0f0f",x"1f1f1f",x"000000",x"000000",
x"0c0c0c",x"1c3971",x"2851a1",x"3060c0",x"224588",x"272727",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"e3e3e3",x"141414",x"000000",x"000000",x"0c1931",x"142951",x"0c1931",x"03060c",
x"2e2e2e",x"8a8a8a",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"e7e7e7",x"dadada",x"ffffff",x"cecece",x"ffffff",x"ffffff",x"cecece",x"bebebe",
x"6e6e6e",x"0e0e0e",x"000000",x"060d19",x"1a1d23",x"d7d7d7",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"cacaca",x"8d8d8d",x"7d7d7d",x"4d4d4d",x"4d4d4d",x"7d7d7d",x"cdcdcd",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"cdcdcd",x"cdcdcd",x"e6e6e6",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",
x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff",x"ffffff"
);
begin
   address <= unsigned(not y(6 downto 0))&unsigned(x(6 downto 0));

process(clk_pixel)
   begin
      if rising_edge(clk_pixel) then
         if a_blank = '0' and pixel /= x"FFFFFF" and x(10 downto 7) = "0000" and y(10 downto 7) = "0000" then
            o_red     <= pixel(7 downto 0);
            o_green   <= pixel(15 downto 8);
            o_blue    <= pixel(23 downto 16);
         else
            o_red     <= a_red;
            o_green   <= a_green;
            o_blue    <= a_blue;
         end if;
         o_blank   <= a_blank;
         o_hsync   <= a_hsync;
         o_vsync   <= a_vsync;

         a_red     <= i_red;
         a_green   <= i_green;
         a_blue    <= i_blue;
         a_blank   <= i_blank;
         a_hsync   <= i_hsync;
         a_vsync   <= i_vsync;

         pixel <= logo(to_integer(address));

         -- Working out where we are in the screen..
         if i_vsync /= a_vsync then
            y <= (others => '0');
         end if;

         if i_blank = '0' then
            x <= std_logic_vector(unsigned(x) + 1);
         end if;

         -- Start of the blanking interval?
         if a_blank = '0' and i_blank = '1' then
            y <= std_logic_vector(unsigned(y) + 1);
            x <= (others => '0');
         end if;

      end if;
   end process;
end Behavioral;

